--! @title     Device Under Test
--! @file      dut.vhd
--! @author    Romain Beaubois
--! @date      29 Nov 2024
--! @copyright
--! SPDX-FileCopyrightText: © 2024 Romain Beaubois <refbeaubois@yahoo.com>
--! SPDX-License-Identifier: MIT
--!
--! @brief Wrapping Wrapping DMA streams and logic with AXI-Lite driven signals
--! * A dummy spike stream in sent to PL via DMA (AXIS SPK_IN) and stored in a FIFO
--! * One time step is read from FIFO at each time step (generated by ts_tick)
--! * Data goes to the black box mimicking actual logic
--! * Processed data is sent back to PS via DMA (AXIS SPK MON)
--! * User LEDs are routed to have all leds lighten when design operates:
--!     - UF1 lighting when bitstream loaded
--!     - UF2 lighting when core enabled
--! 
--! * Simulating AXI-Lite is a pain (pointless extra code and time)
--! so as it's much easier to wrap it this way for simulation
--! 
--! 
--! @details 
--! > **29 Nov 2024** : file creation (RB)

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;

entity dut is
    generic (
        DWIDTH_GPIO         : integer :=    32;
        DWIDTH_DATA         : integer :=    32;
        DWIDTH_SPK_IN       : integer :=    32;
        DWIDTH_SPK_MON      : integer :=    32;
        AWIDTH_FIFO_SPK_IN  : integer :=    10;
        LAT_RD_CDC_FIFO     : integer :=     2;
        MAX_SPK_PER_TS      : integer :=  1000;
        TIME_STEP_CCY       : integer := 12500
    );
    port (
        -- Clock
        clk_pl   : in std_logic;
        clk_axi  : in std_logic;
        srst_pl  : in std_logic;
        srst_axi : in std_logic;
        ts_tick  : out std_logic;

        -- AXI-Lite Control: from PS
        en_core           : in std_logic;

        -- AXI GPIO: from PS
        en_ps_rd_events   : in std_logic;
        ps_rd_events_size : in std_logic_vector(DWIDTH_GPIO-1 downto 0);
        ps_tx_dma_rdy     : in std_logic;

        -- AXI GPIO: to PS
        pl_wr_events_size : out std_logic_vector(DWIDTH_GPIO-1 downto 0);
        count_fifo_spk_in : out std_logic_vector(AWIDTH_FIFO_SPK_IN-1 downto 0);

        -- Spike stream from PS via DMA
        S_AXIS_SPK_IN_ACLK     : in std_logic;
        S_AXIS_SPK_IN_ARESETN  : in std_logic;
        S_AXIS_SPK_IN_TREADY   : out std_logic;
        S_AXIS_SPK_IN_TDATA    : in std_logic_vector(DWIDTH_SPK_IN-1 downto 0);
        S_AXIS_SPK_IN_TLAST    : in std_logic;
        S_AXIS_SPK_IN_TVALID   : in std_logic;

        -- Spike monitoring to DMA
        M_AXIS_SPK_MON_ACLK     : in std_logic;
        M_AXIS_SPK_MON_ARESETN  : in std_logic;
        M_AXIS_SPK_MON_TVALID   : out std_logic;
        M_AXIS_SPK_MON_TREADY   : in std_logic;
        M_AXIS_SPK_MON_TDATA    : out std_logic_vector(DWIDTH_SPK_MON-1 downto 0);
        M_AXIS_SPK_MON_TLAST    : out std_logic;

        -- Periodic interrupts
        ts_pl_wr_ev_intr        : out std_logic;
        
        -- User LEDs
        uled_uf1 : out std_logic;
        uled_uf2 : out std_logic
    );
end entity dut;

architecture rtl of dut is
    -- ========================
    -- Spike stream fed to logic
    -- ========================
    signal raw_rdy_events : std_logic;
    signal raw_ts_event   : std_logic_vector(DWIDTH_SPK_IN-1 downto 0);
    signal raw_nb_event   : std_logic_vector(DWIDTH_SPK_IN-1 downto 0);
    signal raw_id_event   : std_logic_vector(DWIDTH_SPK_IN-1 downto 0);

    -- ========================
    -- Interfacing with logic
    -- ========================
    signal i_logic_rdy_events : std_logic;
    signal i_logic_ts_event   : std_logic_vector(DWIDTH_DATA-1 downto 0);
    signal i_logic_nb_event   : std_logic_vector(DWIDTH_DATA-1 downto 0);
    signal i_logic_id_event   : std_logic_vector(DWIDTH_DATA-1 downto 0);

    signal o_logic_rdy_events : std_logic;
    signal o_logic_ts_event   : std_logic_vector(DWIDTH_DATA-1 downto 0);
    signal o_logic_nb_event   : std_logic_vector(DWIDTH_DATA-1 downto 0);
    signal o_logic_id_event   : std_logic_vector(DWIDTH_DATA-1 downto 0);

    -- ========================
    -- Spike stream processed by logic
    -- ========================
    signal new_rdy_events : std_logic;
    signal new_ts_event   : std_logic_vector(DWIDTH_SPK_MON-1 downto 0);
    signal new_nb_event   : std_logic_vector(DWIDTH_SPK_MON-1 downto 0);
    signal new_id_event   : std_logic_vector(DWIDTH_SPK_MON-1 downto 0);
begin
    ---------------------------------------------------------------------------------------
    --
    --  ████████ ███████     ████████ ██  ██████ ██   ██ 
    --     ██    ██             ██    ██ ██      ██  ██  
    --     ██    ███████        ██    ██ ██      █████   
    --     ██         ██        ██    ██ ██      ██  ██  
    --     ██    ███████        ██    ██  ██████ ██   ██ 
    --
    -- Generate time steps
    ---------------------------------------------------------------------------------------
    timer_proc : process(clk_pl)
        variable cnt : integer range 0 to TIME_STEP_CCY;
    begin
        if rising_edge(clk_pl) then
            if srst_pl = '1' then
                cnt     := TIME_STEP_CCY;
                ts_tick <= '0';
            else
                if en_core = '1' then
                    if cnt > TIME_STEP_CCY-1 then
                        ts_tick <= '1';
                        cnt     := 0;
                    else
                        ts_tick <= '0';
                        cnt     := cnt + 1;
                    end if;
                else
                    ts_tick <= '0';
                    cnt     := TIME_STEP_CCY;
                end if;
            end if;
        end if;
    end process;

    ---------------------------------------------------------------------------------------
    --
    --   █████  ██   ██ ██ ███████     ███████ ██████  ██   ██     ██ ███    ██ 
    --  ██   ██  ██ ██  ██ ██          ██      ██   ██ ██  ██      ██ ████   ██ 
    --  ███████   ███   ██ ███████     ███████ ██████  █████       ██ ██ ██  ██ 
    --  ██   ██  ██ ██  ██      ██          ██ ██      ██  ██      ██ ██  ██ ██ 
    --  ██   ██ ██   ██ ██ ███████     ███████ ██      ██   ██     ██ ██   ████ 
    --                                                                          
    -- Axi signals for Axi subset spikes
    ---------------------------------------------------------------------------------------
    saxis2nat_dma_spk_inst : entity work.saxis2nat_dma_spk_aer
    generic map (
        DWIDTH              => DWIDTH_SPK_IN,
        AWIDTH_FIFO         => AWIDTH_FIFO_SPK_IN,
        LAT_RD_CDC_FIFO     => LAT_RD_CDC_FIFO,
        MAX_SPK_PER_TS      => MAX_SPK_PER_TS
    )
    port map (
        clk_pl                => clk_pl,
        srst_pl               => srst_pl,
        srst_axi              => srst_axi,
        en_core               => en_core,
        ts_tick               => ts_tick,
        ps_tx_dma_rdy         => ps_tx_dma_rdy,
        count_fifo            => count_fifo_spk_in,

        s_axis_aclk           => S_AXIS_SPK_IN_ACLK,
        s_axis_aresetn        => S_AXIS_SPK_IN_ARESETN,
        s_axis_tready         => S_AXIS_SPK_IN_TREADY,
        s_axis_tdata          => S_AXIS_SPK_IN_TDATA,
        s_axis_tlast          => S_AXIS_SPK_IN_TLAST,
        s_axis_tvalid         => S_AXIS_SPK_IN_TVALID,

        rdy_events            => raw_rdy_events,
        ts_event              => raw_ts_event,
        nb_event              => raw_nb_event,
        id_event              => raw_id_event
    );

    ---------------------------------------------------------------------------------------
    --
    --  ██████  ██       █████   ██████ ██   ██ ██████   ██████  ██   ██ 
    --  ██   ██ ██      ██   ██ ██      ██  ██  ██   ██ ██    ██  ██ ██  
    --  ██████  ██      ███████ ██      █████   ██████  ██    ██   ███   
    --  ██   ██ ██      ██   ██ ██      ██  ██  ██   ██ ██    ██  ██ ██  
    --  ██████  ███████ ██   ██  ██████ ██   ██ ██████   ██████  ██   ██ 
    --
    -- Magix blackbox, i.e. your obscure design
    ---------------------------------------------------------------------------------------
    -- Resize data stream from DMA to logic input
    i_logic_rdy_events <= raw_rdy_events;
    i_logic_ts_event   <= std_logic_vector(resize(unsigned(raw_ts_event), DWIDTH_DATA));
    i_logic_nb_event   <= std_logic_vector(resize(unsigned(raw_nb_event), DWIDTH_DATA));
    i_logic_id_event   <= std_logic_vector(resize(unsigned(raw_id_event), DWIDTH_DATA));

    -- Resize data stream from logic input to DMA
    new_rdy_events <= o_logic_rdy_events;
    new_ts_event   <= std_logic_vector(resize(unsigned(o_logic_ts_event), DWIDTH_SPK_MON));
    new_nb_event   <= std_logic_vector(resize(unsigned(o_logic_nb_event), DWIDTH_SPK_MON));
    new_id_event   <= std_logic_vector(resize(unsigned(o_logic_id_event), DWIDTH_SPK_MON));

    -- Instanciate logic module
    blackbox_inst : entity work.blackbox
    generic map(
        DWIDTH_DATA       => DWIDTH_DATA
    )
    port map(
        clk_pl            => clk_pl,
        srst_pl           => srst_pl,

        raw_rdy_in_events => i_logic_rdy_events,
        raw_ts_event      => i_logic_ts_event,
        raw_nb_event      => i_logic_nb_event,
        raw_id_event      => i_logic_id_event,

        new_rdy_in_events => o_logic_rdy_events,
        new_ts_event      => o_logic_ts_event,
        new_nb_event      => o_logic_nb_event,
        new_id_event      => o_logic_id_event
    );

    ---------------------------------------------------------------------------------------
    --                                                                            
    --   █████  ██   ██ ██ ███████     ███████ ██████  ██   ██     ███    ███  ██████  ███    ██ 
    --  ██   ██  ██ ██  ██ ██          ██      ██   ██ ██  ██      ████  ████ ██    ██ ████   ██ 
    --  ███████   ███   ██ ███████     ███████ ██████  █████       ██ ████ ██ ██    ██ ██ ██  ██ 
    --  ██   ██  ██ ██  ██      ██          ██ ██      ██  ██      ██  ██  ██ ██    ██ ██  ██ ██ 
    --  ██   ██ ██   ██ ██ ███████     ███████ ██      ██   ██     ██      ██  ██████  ██   ████ 
    --                                                                                           
    -- Axi signals for Axi subset spikes
    ---------------------------------------------------------------------------------------
    nat2maxis_dma_spk_aer_inst : entity work.nat2maxis_dma_spk_aer
    generic map(
        MAX_SPK_PER_TS  => MAX_SPK_PER_TS,
        DWIDTH_GPIO     => DWIDTH_GPIO,
        DWIDTH_DMA      => DWIDTH_SPK_MON
    )
    port map(
        clk_pl            => clk_pl,
        clk_axi           => clk_axi,
        srst_pl           => srst_pl,
        srst_axi          => srst_axi,
        rdy_in_events     => new_rdy_events,
        ts_event          => new_ts_event,
        nb_event          => new_nb_event,
        id_event          => new_id_event,
        en_ps_rd_events   => en_ps_rd_events,
        pl_wr_events_size => pl_wr_events_size,
        ps_rd_events_size => ps_rd_events_size,
        m_axis_aclk       => M_AXIS_SPK_MON_ACLK,
        m_axis_aresetn    => M_AXIS_SPK_MON_ARESETN,
        m_axis_tvalid     => M_AXIS_SPK_MON_TVALID,
        m_axis_tready     => M_AXIS_SPK_MON_TREADY,
        m_axis_tdata      => M_AXIS_SPK_MON_TDATA,
        m_axis_tlast      => M_AXIS_SPK_MON_TLAST,
        ts_pl_wr_ev_intr  => ts_pl_wr_ev_intr
    );

    ---------------------------------------------------------------------------------------
    --                                                                                   
    --  ██    ██ ███████ ███████ ██████      ██      ███████ ██████  ███████ 
    --  ██    ██ ██      ██      ██   ██     ██      ██      ██   ██ ██      
    --  ██    ██ ███████ █████   ██████      ██      █████   ██   ██ ███████ 
    --  ██    ██      ██ ██      ██   ██     ██      ██      ██   ██      ██ 
    --   ██████  ███████ ███████ ██   ██     ███████ ███████ ██████  ███████ 
    --                                                                                   
    -- User leds for status
    ---------------------------------------------------------------------------------------
    uled_uf1 <= '1';
    uled_uf2 <= en_core;
end architecture;